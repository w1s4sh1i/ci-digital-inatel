/*
Program: CI Digital 02/2025
Class: Introdução à Verilog  
Class-ID: D112
Advisor: Felipe Rocha 
Advisor-Contact: felipef.rocha@inatel.br
Institute: INATEL - Santa Rita do Sapucaí / MG  
Development: André Bezerra 
Student-Contact: andrefrbezerra@gmail.com
Task-ID: A003
Type: Laboratory
Data: octuber, 17 2025
*/

`timescale 1 ns / 1 ps;

module gate_not (
	input signal,
	output not_logic, not_instance
);
	assign not_logic = ~signal;
	not (not_instance, signal);

endmodule
	
