`timescale 1ns/1ps

module codificador_prio_tb();

    reg [15:0] in;
    wire [3:0] out;

    Codificador_Prioridade PRIORITY_TB(
        .in(in),
        .out(out)
    );

    initial begin
        in = 16'b100000000000000; #10;
        in = 16'b010000000000000; #10;
        in = 16'b001000000000000; #10;
        in = 16'b000100000000000; #10;
        in = 16'b000010000000000; #10;
        in = 16'b000001000000000; #10;
        in = 16'b000000100000000; #10;
        in = 16'b000000010000000; #10;
        in = 16'b000000001000000; #10;
        in = 16'b000000000100000; #10;
        in = 16'b000000000010000; #10;
        in = 16'b000000000001000; #10;
        in = 16'b000000000000100; #10;
        in = 16'b000000000000010; #10;
        in = 16'b000000000000001; #10;
        in = 16'b000000000000000; #10;
        $finish;
    end
    

endmodule